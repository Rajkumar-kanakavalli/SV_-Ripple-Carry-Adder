class packet;


randc bit[3:0]a;
randc bit[3:0] b;
randc bit cin;

bit [3:0] sum;
bit cout;

endclass